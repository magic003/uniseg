module main

import os
import net.http
import regex

fn main() {
	if os.args.len < 2 {
		println('Not enough argument. Read code for more details.')
		exit(1)
	}

	segmentation_type := os.args[1]
	match segmentation_type {
		'grapheme' {
			gen_grapheme_properties()
		}
		else {
			println('Unrecognized argument: ${segmentation_type}')
			exit(1)
		}
	}
}

// unicode_version is the Unicode version that this unicode-segmentation lib is based on.
const unicode_version = '15.0.0'

const (
	grapheme_property_url = 'https://www.unicode.org/Public/${unicode_version}/ucd/auxiliary/GraphemeBreakProperty.txt'
	emoji_property_url    = 'https://unicode.org/Public/${unicode_version}/ucd/emoji/emoji-data.txt'
)

// property_line_regex is the regexp matching a property line.
const property_line_regex = r'^(?P<start>[0-9A-F]{4,6})(\.\.(?P<to>[0-9A-F]{4,6}))?\s*;\s*(?P<property>[A-Za-z0-9_]+)\s*#\s(?P<comment>.+)$'

// Property represents a property. It is a line in the fetched properties file.
struct Property {
	from    string
	to      string
	name    string
	comment string
}

fn gen_grapheme_properties() {
	mut properties := []Property{}

	properties << parse_properties(grapheme_property_url, fn (line string) bool {
		return true
	})

	properties << parse_properties(emoji_property_url, fn (line string) bool {
		return line.contains('Extended_Pictographic')
	})

	properties.sort(a.from < b.from)

	write_grapheme_properties(properties) or { panic(error) }
}

fn parse_properties(url string, filter fn (string) bool) []Property {
	mut properties := []Property{}

	println('Fetching ${url}...')
	lines := http.get_text(url).split_into_lines()
	for line in lines {
		if line.len == 0 || line.starts_with('#') || !filter(line) {
			continue
		}
		prop := parse_line(line) or { continue }
		properties << prop
	}
	println('Finish parsing ${url}.')

	return properties
}

fn parse_line(line string) ?Property {
	mut re := regex.regex_opt(property_line_regex) or { panic(error) }
	match_start, _ := re.match_string(line)
	if match_start < 0 {
		return none
	}

	from := re.get_group_by_name(line, 'start')
	to_group := re.get_group_by_name(line, 'to')
	to := if to_group != '' {
		to_group
	} else {
		from
	}
	property := re.get_group_by_name(line, 'property')
	comment := re.get_group_by_name(line, 'comment')

	return Property{from, to, property, comment}
}

fn write_grapheme_properties(properties []Property) ! {
	vfile_path := 'src/grapheme/grapheme_properties.v'
	println('Saving to file ${vfile_path}...')
	mut file := os.create(vfile_path)!
	defer {
		file.close()
		println('Finish saving file ${vfile_path}.')
	}
	file.writeln(emit_module('grapheme') + '\n')!
	file.writeln(emit_preamble() + '\n')!
	file.writeln(emit_property_enum('GraphemeProp', unique_property_names(properties), 'gp') + '\n')!
	file.writeln(emit_code_points_struct('GraphemeCodePoint', 'GraphemeProp') + '\n')!
	file.writeln(emit_property_array(properties, 'GraphemeCodePoint', 'GraphemeProp', 'gp') + '\n')!
}

fn unique_property_names(properties []Property) []string {
	mut res := []string{}
	mut prop_set := map[string]Property{}
	for prop in properties {
		if prop.name !in prop_set {
			prop_set[prop.name] = prop
			res << prop.name
		}
	}

	return res
}

fn emit_module(mod string) string {
	return 'module ${mod}'
}

fn emit_preamble() string {
	return '// NOTE: The following code was generated by "gen/gen_properties.v". DO NOT EDIT.'
}

fn emit_property_enum(name string, values []string, prefix string) string {
	mut res := 'enum ${name} {\n'
	res += '\t${prefix}_any\n'
	for v in values {
		res += '\t${prefix}_${v.to_lower()}\n'
	}
	res += '}'

	return res
}

fn emit_code_points_struct(name string, property_enum_name string) string {
	mut res := 'struct ${name} {\n'
	res += '\tfrom int\n'
	res += '\tto int\n'
	res += '\tproperty ${property_enum_name}\n'
	res += '}'
	return res
}

fn emit_property_array(properties []Property, code_point_struct_name string, enum_name string, prefix string) string {
	mut res := 'const grapheme_properties = [\n'
	for prop in properties {
		res += '\t${code_point_struct_name}{0x${prop.from}, 0x${prop.to}, ${enum_name}.${prefix}_${prop.name.to_lower()}},\n'
	}
	res += ']'
	return res
}
