module common

import datatypes
import net.http
import regex

// unicode_version is the Unicode version that this unicode-segmentation lib is based on.
pub const unicode_version = '15.0.0'

// property_line_regex is the regexp matching a property line.
const property_line_regex = r'^(?P<start>[0-9A-F]{4,6})(\.\.(?P<to>[0-9A-F]{4,6}))?\s*;\s*(?P<property>[A-Za-z0-9_]+)\s*#\s(?P<comment>.+)$'

// Property represents a property. It is a line in the fetched properties file.
pub struct Property {
pub:
	from    string
	to      string
	name    string
	comment string
}

// parse_properties parses the property file in a URL into an array of properties.
pub fn parse_properties(url string, filter fn (string) bool) []Property {
	mut properties := []Property{}

	println('Fetching ${url}...')
	lines := http.get_text(url).split_into_lines()
	for line in lines {
		if line.len == 0 || line.starts_with('#') || !filter(line) {
			continue
		}
		prop := parse_line(line) or { continue }
		properties << prop
	}
	println('Finish parsing ${url}.')

	return properties
}

// parse_line parses a single line in a property file.
fn parse_line(line string) ?Property {
	mut re := regex.regex_opt(common.property_line_regex) or { panic(error) }
	match_start, _ := re.match_string(line)
	if match_start < 0 {
		return none
	}

	from := re.get_group_by_name(line, 'start')
	to_group := re.get_group_by_name(line, 'to')
	to := if to_group != '' {
		to_group
	} else {
		from
	}
	property := re.get_group_by_name(line, 'property')
	comment := re.get_group_by_name(line, 'comment')

	return Property{from, to, property, comment}
}

// unique_property_names extract the unique names from an array of properties, in the same order.
pub fn unique_property_names(properties []Property) []string {
	mut res := []string{}
	mut prop_set := datatypes.Set[string]{}
	for prop in properties {
		if !prop_set.exists(prop.name) {
			prop_set.add(prop.name)
			res << prop.name
		}
	}

	return res
}

// emit_module generates a vlang module statement.
pub fn emit_module(mod string) string {
	return 'module ${mod}'
}

// emit_preamble generates a preamble for a vlang file.
pub fn emit_preamble(script string) string {
	return '// NOTE: The following code was generated by "${script}". DO NOT EDIT.'
}

// emit_property_enum generates a vlang `enum` for property types.
pub fn emit_property_enum(name string, values []string, prefix string) string {
	mut res := 'enum ${name} {\n'
	res += '\t${prefix}_any\n'
	for v in values {
		res += '\t${prefix}_${v.to_lower()}\n'
	}
	res += '}'

	return res
}

// emit_code_points_struct generates a vlang `struct` for code points.
pub fn emit_code_points_struct(name string, property_enum_name string) string {
	mut res := 'struct ${name} {\n'
	res += '\tfrom int\n'
	res += '\tto int\n'
	res += '\tproperty ${property_enum_name}\n'
	res += '}'
	return res
}

// emit_property_array generates a vlang `array` of particular properties.
pub fn emit_property_array(name string, properties []Property, code_point_struct_name string, enum_name string, prefix string) string {
	mut res := 'const ${name} = [\n'
	for prop in properties {
		res += '\t${code_point_struct_name}{0x${prop.from}, 0x${prop.to}, ${enum_name}.${prefix}_${prop.name.to_lower()}}, // ${prop.comment}\n'
	}
	res += ']'
	return res
}
